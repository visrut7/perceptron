module matrix

pub type Matrix = [][]f64
